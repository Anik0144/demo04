magic
tech sky130A
timestamp 1680899189
<< nwell >>
rect -70 135 85 335
<< pwell >>
rect -95 -40 110 100
<< nmos >>
rect 0 -30 15 70
<< pmos >>
rect 0 155 15 309
<< ndiff >>
rect -40 55 0 70
rect -40 -15 -35 55
rect -15 -15 0 55
rect -40 -30 0 -15
rect 15 55 55 70
rect 15 -15 30 55
rect 50 -15 55 55
rect 15 -30 55 -15
<< pdiff >>
rect -45 290 0 309
rect -45 170 -35 290
rect -15 170 0 290
rect -45 155 0 170
rect 15 290 60 309
rect 15 175 30 290
rect 50 175 60 290
rect 15 155 60 175
<< ndiffc >>
rect -35 -15 -15 55
rect 30 -15 50 55
<< pdiffc >>
rect -35 170 -15 290
rect 30 175 50 290
<< poly >>
rect 0 309 15 395
rect 0 125 15 155
rect -45 115 15 125
rect -45 90 -35 115
rect -5 90 15 115
rect -45 80 15 90
rect 0 70 15 80
rect 0 -55 15 -30
<< polycont >>
rect -35 90 -5 115
<< locali >>
rect -40 482 85 496
rect -40 436 -28 482
rect 67 436 85 482
rect -40 426 85 436
rect -35 290 -15 426
rect -35 155 -15 170
rect 30 300 50 305
rect 30 290 55 300
rect 50 175 55 290
rect 30 135 55 175
rect -55 90 -35 115
rect -5 90 15 115
rect 35 70 55 135
rect -35 55 -15 70
rect -35 -85 -15 -15
rect 30 55 55 70
rect 50 -15 55 55
rect 30 -30 55 -15
rect -50 -95 70 -85
rect -50 -120 -40 -95
rect 60 -120 70 -95
rect -50 -130 70 -120
<< viali >>
rect -28 436 67 482
rect -40 -120 60 -95
<< metal1 >>
rect -51 482 93 500
rect -51 436 -28 482
rect 67 436 93 482
rect -51 425 93 436
rect -50 -95 70 -85
rect -50 -120 -40 -95
rect 60 -120 70 -95
rect -50 -130 70 -120
<< end >>
