magic
tech sky130A
timestamp 1675131467
<< error_p >>
rect -3 145 5 153
rect 8 137 13 145
rect 8 133 10 137
rect 8 125 13 133
rect -3 117 5 125
rect 25 108 27 162
<< nwell >>
rect -70 150 80 365
<< pwell >>
rect -70 115 85 120
rect -70 110 -25 115
rect 0 110 85 115
rect -70 -30 85 110
<< nmos >>
rect 0 0 15 100
<< pmos >>
rect 0 170 15 346
<< ndiff >>
rect -40 90 0 100
rect -40 5 -30 90
rect -10 5 0 90
rect -40 0 0 5
rect 15 95 55 100
rect 15 5 25 95
rect 45 5 55 95
rect 15 0 55 5
<< pdiff >>
rect -35 335 0 346
rect -35 180 -30 335
rect -10 180 0 335
rect -35 170 0 180
rect 15 335 50 346
rect 15 180 25 335
rect 45 180 50 335
rect 15 170 50 180
<< ndiffc >>
rect -30 5 -10 90
rect 25 5 45 95
<< pdiffc >>
rect -30 180 -10 335
rect 25 180 45 335
<< poly >>
rect 0 346 15 375
rect 0 155 15 170
rect -30 145 15 155
rect -30 125 -25 145
rect 5 125 15 145
rect -30 115 15 125
rect 0 100 15 115
rect 0 -20 15 0
<< polycont >>
rect -25 125 5 145
<< locali >>
rect -80 370 95 405
rect -30 335 -10 370
rect -30 170 -10 180
rect 25 335 45 345
rect 25 175 45 180
rect -35 125 -25 145
rect 5 125 10 145
rect 25 100 60 175
rect -30 90 -10 100
rect -30 -30 -10 5
rect 25 95 45 100
rect 25 -5 45 5
rect -70 -70 85 -30
<< end >>
